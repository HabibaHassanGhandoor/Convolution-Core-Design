`timescale 1ns/1ns

module top_tb;

  // Define constants
  parameter CLK_PERIOD = 10; // Clock period in ns

  // Declare signals for the testbench
  reg clk, rst;
  reg [127:0] Datain;
  reg [1:0] control;
  wire Valid, Done;
  wire [127:0] Dataout;
  wire invalid_operation;

  // Instantiate the top module
  top uut (
    .clk(clk),
    .rst(rst),
    .Datain(Datain),
    .control(control),
    .Valid(Valid),
    .Done(Done),
    .Dataout(Dataout),
    .invalid_operation(invalid_operation)
  );

  // Clock generation
  always begin
    #(CLK_PERIOD/2) clk = ~clk; // Toggle the clock
  end

  // Initial block for simulation setup
  initial begin
    // Initialize signals
    clk = 0;
    rst = 0; // Active-low reset

    // Apply reset for a few clock cycles
    #20 rst = 1;
    //test case 1 no floating point or negative
    //load configurations
    //input matrix 3*3   kernel matrix 2*2     stride=1
    Datain[7:0] = 8'd2;   //M
		Datain[15:8] = 8'd2;  //N
		Datain[23:16] = 8'd1;  //S
		Datain[31:24] = 8'd3;  //L
		Datain[39:32] = 8'd3;  //W
	  Datain [127:40] = 'b0;
	  control = 2'b00; // Set initial value for control
	  #50
	  
	  
	  //load kernel
	  Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
    control = 2'b01;
    #10;
  
    
    //load input
    control = 2'b10; 
    Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  
 #10
	  Datain[31:0] = 32'b01000000100000000000000000000000;  //4
	  Datain[63:32] = 32'b01000000101000000000000000000000;  //5
	  Datain[95:64] = 32'b01000000110000000000000000000000;  //6
	  Datain [127:96] = 32'b01000000111000000000000000000000; //7
	  #10
	  Datain[31:0] = 32'b01000001000000000000000000000000;  //8
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  #10
	  control = 2'b11;
	  
    #400
    
    ///testing remaider = 1
    
        //load configurations
    //input matrix 3*3   kernel matrix 2*2     stride=2
    Datain[7:0] = 8'd2;   //M
		Datain[15:8] = 8'd2;  //N
		Datain[23:16] = 8'd2;  //S
		Datain[31:24] = 8'd3;  //L
		Datain[39:32] = 8'd3;  //W
	  Datain [127:40] = 'b0;
	  control = 2'b00; // Set initial value for control
	  #50
	  
	  
	  //load kernel
	  Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
    control = 2'b01;
    #10;
  
    
    //load input
    control = 2'b10; 
    Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  
 #10
	  Datain[31:0] = 32'b01000000100000000000000000000000;  //4
	  Datain[63:32] = 32'b01000000101000000000000000000000;  //5
	  Datain[95:64] = 32'b01000000110000000000000000000000;  //6
	  Datain [127:96] = 32'b01000000111000000000000000000000; //7
	  #10
	  Datain[31:0] = 32'b01000001000000000000000000000000;  //8
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  #10
	  control = 2'b11;
				
    #400
    
    ///testing kernel with  negative values and input with floating point values
    
        //load configurations
    //input matrix 5*5   kernel matrix 3*3     stride=1
    Datain[7:0] = 8'd3;   //M
		Datain[15:8] = 8'd3;  //N
		Datain[23:16] = 8'd1;  //S
		Datain[31:24] = 8'd5;  //L
		Datain[39:32] = 8'd5;  //W
	  Datain [127:40] = 'b0;
	  control = 2'b00; // Set initial value for control
	  #50
	  
	  
	  //load kernel
	  Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b10111111100000000000000000000000;  //-1
	  Datain[95:64] = 32'b00000000000000000000000000000000;  //0
	  Datain [127:96] = 32'b10111111100000000000000000000000; //-1
    control = 2'b01;
    #10;
    Datain[31:0] = 32'b01000000101000000000000000000000;  //5
	  Datain[63:32] = 32'b10111111100000000000000000000000;  //-1
	  Datain[95:64] = 32'b00000000000000000000000000000000;  //0
	  Datain [127:96] = 32'b10111111100000000000000000000000; //-1
    #10;
    Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b10111111100000000000000000000000;  //-1
	  Datain[95:64] = 32'b00000000000000000000000000000000;  //0
	  Datain [127:96] = 32'b10111111100000000000000000000000; //-1
    #10
  
    
    //load input
    control = 2'b10; 
    Datain[31:0] = 32'b00111110010011001100110011001101;  //0.2
	  Datain[63:32] = 32'b00111110110011001100110011001101;  //0.4
	  Datain[95:64] = 32'b00111111000110011001100110011010;  //0.6
	  Datain [127:96] = 32'b00111111010011001100110011001101; //0.8
	  
    #10
	  Datain[31:0] = 32'b00111111100000000000000000000000;  //1
	  Datain[63:32] = 32'b00111101110011001100110011001101;  //0.1
	  Datain[95:64] = 32'b00111110100110011001100110011010;  //0.3                 
	  Datain [127:96] = 32'b00111111000000000000000000000000; //0.5
	  #10
	  Datain[31:0] = 32'b00111111001100110011001100110011;  //0.7
	  Datain[63:32] = 32'b00111111011001100110011001100110;  //0.9
	  Datain[95:64] = 32'b00000000000000000000000000000000;  //0
	  Datain [127:96] = 32'b00111110010011001100110011001101; //0.2  
	  #10
	  Datain[31:0] = 32'b00111110110011001100110011001101;  //0.4
	  Datain[63:32] = 32'b00111111000110011001100110011010;  //0.6
	  Datain [95:64] = 32'b00111111010011001100110011001101; //0.8
	  Datain [127:96] = 32'b00111101110011001100110011001101; //0.1
	  #10
	  Datain[31:0] = 32'b00111110100110011001100110011010;  //0.3
	  Datain[63:32] = 32'b00111111000000000000000000000000;  //0.5
	  Datain [95:64] = 32'b00111111001100110011001100110011; //0.7
	  Datain [127:96] = 32'b00111111011001100110011001100110; //0.9
	  #10
	  Datain[31:0] = 32'b00111110010011001100110011001101;  //0.2
	  Datain[63:32] = 32'b00111110110011001100110011001101;  //0.4
	  Datain[95:64] = 32'b00111111000110011001100110011010;  //0.6
	  Datain [127:96] = 32'b00111111010011001100110011001101; //0.8
    #10
    Datain[31:0] = 32'b00111111100000000000000000000000;  //1
	  Datain[63:32] = 32'b00111101110011001100110011001101;  //0.1
	  Datain[95:64] = 32'b00111110100110011001100110011010;  //0.3
	  Datain [127:96] = 32'b00111111000000000000000000000000; //0.5
	  #10
    
	  
	  control = 2'b11;
				
    #1000
    
//    //testing invalid_operation signal (not square matrix)
//    Datain[7:0] = 8'd2;   //M
//		Datain[15:8] = 8'd2;  //N
//		Datain[23:16] = 8'd1;  //S
//		Datain[31:24] = 8'd3;  //L
//		Datain[39:32] = 8'd2;  //W
//	  Datain [127:40] = 'b0;
//	  control = 2'b00; // Set initial value for control
//	  #50
//	  //load kernel
//	  Datain[31:0] = 32'b00000000000000000000000000000000;  //0
//	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
//	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
//	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
//    control = 2'b01;
//    #10;
//  
//    
//    //load input
//    control = 2'b10; 
//    Datain[31:0] = 32'b00000000000000000000000000000000;  //0
//	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
//	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
//	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
//	  
//    #10
//	  Datain[31:0] = 32'b01000000100000000000000000000000;  //4
//	  Datain[63:32] = 32'b01000000101000000000000000000000;  //5
//	  Datain[95:64] = 32'b01000000110000000000000000000000;  //6
//	  Datain [127:96] = 32'b01000000111000000000000000000000; //7
//	  #10
//
//	  control = 2'b11;
//	  
//    #400
    
    //testing invalid_operation signal (kernel size is larger than input size)
    Datain[7:0] = 8'd3;   //M
		Datain[15:8] = 8'd3;  //N
		Datain[23:16] = 8'd1;  //S
		Datain[31:24] = 8'd2;  //L
		Datain[39:32] = 8'd2;  //W
	  Datain [127:40] = 'b0;
	  control = 2'b00; // Set initial value for control
	  #50
	  //load kernel
	  Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
    control = 2'b01;
    #10
	  Datain[31:0] = 32'b01000000100000000000000000000000;  //4
	  Datain[63:32] = 32'b01000000101000000000000000000000;  //5
	  Datain[95:64] = 32'b01000000110000000000000000000000;  //6
	  Datain [127:96] = 32'b01000000111000000000000000000000; //7
    #10
	  Datain[31:0] = 32'b01000001000000000000000000000000;  //8
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  #10
  
    
    //load input
    control = 2'b10; 
    Datain[31:0] = 32'b00000000000000000000000000000000;  //0
	  Datain[63:32] = 32'b00111111100000000000000000000000;  //1
	  Datain[95:64] = 32'b01000000000000000000000000000000;  //2
	  Datain [127:96] = 32'b01000000010000000000000000000000; //3
	  
	  #10

	  control = 2'b11;
	  
    #400
    
    
    $stop; // Stop the simulation after 1000 time units

  end

endmodule



